module adder (
    ports
);
    
endmodule